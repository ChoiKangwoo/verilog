/*It is a 4-bit parallel adder module using a 4 bit carry-lookahead module*/
module AdderCLA(a,b,cin,sum,cout);


//Input declaration

	//Declare array a,b with size 4
	input [3:0] a,b;

	//c0=cin
	input cin;

//Output declaration

	//Declare array sum with size 4	
	output [3:0] sum;

	//c4=cout
	output cout;

//wire declaration

	//Array with a size of 4 that stores the Carry value
	wire [4:1] C;

	//Declare an array with a size of 4 storing G,P
	wire [3:0] G;
	wire [3:0] P;

//FullAdder Operation Interval

	//First bit calculation, G0 and P0 are output.
	fulladder A1 (a[0],b[0],cin,sum[0],G[0],P[0]);

	//Second bit calculation, G1 and P1 are output.
	fulladder A2 (a[1],b[1],C[1],sum[1],G[1],P[1]);

	//Third bit calculation, G2 and P2 are output.
	fulladder A3 (a[2],b[2],C[2],sum[2],G[2],P[2]);

	//Fourth bit calculation, G3 and P3 are output.
	fulladder A4 (a[3],b[3],C[3],sum[3],G[3],P[3]);

//CLA Operation Interval

	//G0, G1, G2, G3 and P0, P1, P2, and P3 calculated by the adder are received 
	//and C1, C2, C3, and C4 are output.
	//cin is c0
	CLA C1 (G,P,cin,C);

	assign cout= C[4];

	
	
	
	


endmodule

/*It is an adder module that outputs G and P values and 
calculates the sum.*/

module fulladder(a,b,cin,sum,Gout,Pout);

	input a,b,cin;

	output sum;
	output Gout,Pout;
	
	//calculates the sum with operated by XOR gate.
	assign sum=a^b^cin;
	
	//Gi=Ai&Bi ; indicates the ith stage generate a carryout
	assign Gout=a&b;

	//Pi=Ai^Bi ; indicates the ith stage propagate a carry into carryout
	assign Pout=a^b;

endmodule


/*By receiving the calculated G and P values, 
the carrier values generated by the addition of A and B are calculated.
 */
module CLA (G,P,cin,cout);
	

	input [3:0] G,P;
	input cin;
	
	output [4:1] cout;
	

	//calculate using carry-lookahead equation 
	assign cout[1]=G[0] | P[0]&cin;
	assign cout[2]=G[1] | P[1]&G[0]| P[1]&P[0]&cin;
	assign cout[3]=G[2] | P[2]&G[1]| P[2]&P[1]&G[0]| P[2]&P[1]&P[0]&cin;
	assign cout[4]=G[3] | P[3]&G[2] | P[3]&P[2]&G[1]|P[3]&P[2]&P[1]&G[0]|P[3]&P[2]&P[1]&P[0]&cin;
endmodule






